// Automatically generated Verilog-2001
module MatrixMultiplyCore3x3_busBuild14(ds
                                       ,result);
  input [19:0] ds;
  output [19:0] result;
  assign result = ds + 20'd1;
endmodule
