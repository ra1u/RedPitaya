// Automatically generated Verilog-2001
module MatrixMultiplyCore3x3_BitPackBitVector1(v
                                              ,result);
  input [0:0] v;
  output [0:0] result;
  assign result = v;
endmodule
